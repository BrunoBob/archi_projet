--ALU
